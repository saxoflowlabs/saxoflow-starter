Formal property generation commented out.